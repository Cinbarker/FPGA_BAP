library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity project_toplevel is
--  Port ( );
end project_toplevel;

architecture behavioral of project_toplevel is

begin


end behavioral;
